`include "timescale.v"
module tst_bench_top(); reg clk; reg rstn; wire [31:0] adr; wire [ 7:0] dat_i, dat_o, dat0_i, dat1_i; wire we; wire stb; wire cyc; wire ack; wire inta; reg [7:0] q, qq; wire scl, scl0_o, scl0_oen, scl1_o, scl1_oen; wire sda, sda0_o, sda0_oen, sda1_o, sda1_oen; parameter PRER_LO = 3'b000; parameter PRER_HI = 3'b001; parameter CTR = 3'b010; parameter RXR = 3'b011; parameter TXR = 3'b011; parameter CR = 3'b100; parameter SR = 3'b100; parameter TXR_R = 3'b101; parameter CR_R = 3'b110; parameter RD = 1'b1; parameter WR = 1'b0; parameter SADR = 7'b0010_000; always #5 clk = ~clk; wb_master_model #(8, 32) u0 ( .clk(clk), .rst(rstn), .adr(adr), .din(dat_i), .dout(dat_o), .cyc(cyc), .stb(stb), .we(we), .sel(), .ack(ack), .err(1'b0), .rty(1'b0) ); wire stb0 = stb & ~adr[3]; wire stb1 = stb & adr[3]; assign dat_i = ({{8'd8}{stb0}} & dat0_i) | ({{8'd8}{stb1}} & dat1_i); i2c_master_top i2c_top ( .wb_clk_i(clk), .wb_rst_i(1'b0), .arst_i(rstn), .wb_adr_i(adr[2:0]), .wb_dat_i(dat_o), .wb_dat_o(dat0_i), .wb_we_i(we), .wb_stb_i(stb0), .wb_cyc_i(cyc), .wb_ack_o(ack), .wb_inta_o(inta), .scl_pad_i(scl), .scl_pad_o(scl0_o), .scl_padoen_o(scl0_oen), .sda_pad_i(sda), .sda_pad_o(sda0_o), .sda_padoen_o(sda0_oen) ), i2c_top2 ( .wb_clk_i(clk), .wb_rst_i(1'b0), .arst_i(rstn), .wb_adr_i(adr[2:0]), .wb_dat_i(dat_o), .wb_dat_o(dat1_i), .wb_we_i(we), .wb_stb_i(stb1), .wb_cyc_i(cyc), .wb_ack_o(ack), .wb_inta_o(inta), .scl_pad_i(scl), .scl_pad_o(scl1_o), .scl_padoen_o(scl1_oen), .sda_pad_i(sda), .sda_pad_o(sda1_o), .sda_padoen_o(sda1_oen) ); i2c_slave_model #(SADR) i2c_slave ( .scl(scl), .sda(sda) ); delay m0_scl (scl0_oen ? 1'bz : scl0_o, scl), m1_scl (scl1_oen ? 1'bz : scl1_o, scl), m0_sda (sda0_oen ? 1'bz : sda0_o, sda), m1_sda (sda1_oen ? 1'bz : sda1_o, sda); pullup p1(scl); pullup p2(sda); initial begin `ifdef WAVES
$shm_open("waves"); $shm_probe("AS",tst_bench_top,"AS"); $display("INFO: Signal dump enabled ...\n\n"); `endif
force i2c_slave.debug = 1'b0; $display("\nstatus: %t Testbench started\n\n", $time); clk = 0; rstn = 1'b1; #2; rstn = 1'b0; repeat(1) @(posedge clk); rstn = 1'b1; $display("status: %t done reset", $time); @(posedge clk); u0.wb_write(1, PRER_LO, 8'hfa); u0.wb_write(1, PRER_LO, 8'hc8); u0.wb_write(1, PRER_HI, 8'h00); $display("status: %t programmed registers", $time); u0.wb_cmp(0, PRER_LO, 8'hc8); u0.wb_cmp(0, PRER_HI, 8'h00); $display("status: %t verified registers", $time); u0.wb_write(1, CTR, 8'h80); $display("status: %t core enabled", $time); u0.wb_write(1, TXR, {SADR,WR} ); u0.wb_write(0, CR, 8'h90 ); $display("status: %t generate 'start', write cmd %0h (slave address+write)", $time, {SADR,WR} ); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(0, SR, q); $display("status: %t tip==0", $time); u0.wb_write(1, TXR, 8'h01); u0.wb_write(0, CR, 8'h10); $display("status: %t write slave memory address 01", $time); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(0, SR, q); $display("status: %t tip==0", $time); u0.wb_write(1, TXR, 8'ha5); u0.wb_write(0, CR, 8'h10); $display("status: %t write data a5", $time); while (scl) #1; force scl= 1'b0; #100000; release scl; u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_write(1, TXR, 8'h5a); u0.wb_write(0, CR, 8'h50); $display("status: %t write next data 5a, generate 'stop'", $time); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_write(1, TXR,{SADR,WR} ); u0.wb_write(0, CR, 8'h90 ); $display("status: %t generate 'start', write cmd %0h (slave address+write)", $time, {SADR,WR} ); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_write(1, TXR, 8'h01); u0.wb_write(0, CR, 8'h10); $display("status: %t write slave address 01", $time); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_write(1, TXR, {SADR,RD} ); u0.wb_write(0, CR, 8'h90 ); $display("status: %t generate 'repeated start', write cmd %0h (slave address+read)", $time, {SADR,RD} ); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_write(1, CR, 8'h20); $display("status: %t read + ack", $time); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_read(1, RXR, qq); if(qq !== 8'ha5) $display("\nERROR: Expected a5, received %x at time %t", qq, $time); else $display("status: %t received %x", $time, qq); u0.wb_write(1, CR, 8'h20); $display("status: %t read + ack", $time); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_read(1, RXR, qq); if(qq !== 8'h5a) $display("\nERROR: Expected 5a, received %x at time %t", qq, $time); else $display("status: %t received %x", $time, qq); u0.wb_write(1, CR, 8'h20); $display("status: %t read + ack", $time); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_read(1, RXR, qq); $display("status: %t received %x from 3rd read address", $time, qq); u0.wb_write(1, CR, 8'h28); $display("status: %t read + nack", $time); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_read(1, RXR, qq); $display("status: %t received %x from 4th read address", $time, qq); u0.wb_write(1, TXR, {SADR,WR} ); u0.wb_write(0, CR, 8'h90 ); $display("status: %t generate 'start', write cmd %0h (slave address+write). Check invalid address", $time, {SADR,WR} ); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); u0.wb_write(1, TXR, 8'h10); u0.wb_write(0, CR, 8'h10); $display("status: %t write slave memory address 10", $time); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); $display("status: %t Check for nack", $time); if(!q[7]) $display("\nERROR: Expected NACK, received ACK\n"); u0.wb_write(1, CR, 8'h40); $display("status: %t generate 'stop'", $time); u0.wb_read(1, SR, q); while(q[1]) u0.wb_read(1, SR, q); $display("status: %t tip==0", $time); #250000; $display("\n\nstatus: %t Testbench done", $time); $finish; end endmodule module delay (in, out); input in; output out; assign out = in; specify (in => out) = (600,600); endspecify endmodule