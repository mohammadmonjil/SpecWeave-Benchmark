// Auto-flattened Verilog file

// ===== Macros =====
`define I2C_CMD_NOP 4'b0000
`define I2C_CMD_START 4'b0001
`define I2C_CMD_STOP 4'b0010
`define I2C_CMD_WRITE 4'b0100
`define I2C_CMD_READ 4'b1000


// ==== Module: i2c_master_top ====
module i2c_master_top( wb_clk_i, wb_rst_i, arst_i, wb_adr_i, wb_dat_i, wb_dat_o, wb_we_i, wb_stb_i, wb_cyc_i, wb_ack_o, wb_inta_o, scl_pad_i, scl_pad_o, scl_padoen_o, sda_pad_i, sda_pad_o, sda_padoen_o ); parameter ARST_LVL = 1'b0; input wb_clk_i; input wb_rst_i; input arst_i; input [2:0] wb_adr_i; input [7:0] wb_dat_i; output [7:0] wb_dat_o; input wb_we_i; input wb_stb_i; input wb_cyc_i; output wb_ack_o; output wb_inta_o; reg [7:0] wb_dat_o; reg wb_ack_o; reg wb_inta_o; input scl_pad_i; output scl_pad_o; output scl_padoen_o; input sda_pad_i; output sda_pad_o; output sda_padoen_o; reg [15:0] prer; reg [ 7:0] ctr; reg [ 7:0] txr; wire [ 7:0] rxr; reg [ 7:0] cr; wire [ 7:0] sr; wire done; wire core_en; wire ien; wire irxack; reg rxack; reg tip; reg irq_flag; wire i2c_busy; wire i2c_al; reg al; wire rst_i = arst_i ^ ARST_LVL; wire wb_wacc = wb_we_i & wb_ack_o; always @(posedge wb_clk_i) wb_ack_o <= #1 wb_cyc_i & wb_stb_i & ~wb_ack_o; always @(posedge wb_clk_i) begin case (wb_adr_i) 3'b000: wb_dat_o <= #1 prer[ 7:0]; 3'b001: wb_dat_o <= #1 prer[15:8]; 3'b010: wb_dat_o <= #1 ctr; 3'b011: wb_dat_o <= #1 rxr; 3'b100: wb_dat_o <= #1 sr; 3'b101: wb_dat_o <= #1 txr; 3'b110: wb_dat_o <= #1 cr; 3'b111: wb_dat_o <= #1 0; endcase end always @(posedge wb_clk_i or negedge rst_i) if (!rst_i) begin prer <= #1 16'hffff; ctr <= #1 8'h0; txr <= #1 8'h0; end else if (wb_rst_i) begin prer <= #1 16'hffff; ctr <= #1 8'h0; txr <= #1 8'h0; end else if (wb_wacc) case (wb_adr_i) 3'b000 : prer [ 7:0] <= #1 wb_dat_i; 3'b001 : prer [15:8] <= #1 wb_dat_i; 3'b010 : ctr <= #1 wb_dat_i; 3'b011 : txr <= #1 wb_dat_i; default: ; endcase always @(posedge wb_clk_i or negedge rst_i) if (!rst_i) cr <= #1 8'h0; else if (wb_rst_i) cr <= #1 8'h0; else if (wb_wacc) begin if (core_en & (wb_adr_i == 3'b100) ) cr <= #1 wb_dat_i; end else begin if (done | i2c_al) cr[7:4] <= #1 4'h0; cr[2:1] <= #1 2'b0; cr[0] <= #1 1'b0; end wire sta = cr[7]; wire sto = cr[6]; wire rd = cr[5]; wire wr = cr[4]; wire ack = cr[3]; wire iack = cr[0]; assign core_en = ctr[7]; assign ien = ctr[6]; i2c_master_byte_ctrl byte_controller ( .clk ( wb_clk_i ), .rst ( wb_rst_i ), .nReset ( rst_i ), .ena ( core_en ), .clk_cnt ( prer ), .start ( sta ), .stop ( sto ), .read ( rd ), .write ( wr ), .ack_in ( ack ), .din ( txr ), .cmd_ack ( done ), .ack_out ( irxack ), .dout ( rxr ), .i2c_busy ( i2c_busy ), .i2c_al ( i2c_al ), .scl_i ( scl_pad_i ), .scl_o ( scl_pad_o ), .scl_oen ( scl_padoen_o ), .sda_i ( sda_pad_i ), .sda_o ( sda_pad_o ), .sda_oen ( sda_padoen_o ) ); always @(posedge wb_clk_i or negedge rst_i) if (!rst_i) begin al <= #1 1'b0; rxack <= #1 1'b0; tip <= #1 1'b0; irq_flag <= #1 1'b0; end else if (wb_rst_i) begin al <= #1 1'b0; rxack <= #1 1'b0; tip <= #1 1'b0; irq_flag <= #1 1'b0; end else begin al <= #1 i2c_al | (al & ~sta); rxack <= #1 irxack; tip <= #1 (rd | wr); irq_flag <= #1 (done | i2c_al | irq_flag) & ~iack; end always @(posedge wb_clk_i or negedge rst_i) if (!rst_i) wb_inta_o <= #1 1'b0; else if (wb_rst_i) wb_inta_o <= #1 1'b0; else wb_inta_o <= #1 irq_flag && ien; assign sr[7] = rxack; assign sr[6] = i2c_busy; assign sr[5] = al; assign sr[4:2] = 3'h0; assign sr[1] = tip; assign sr[0] = irq_flag; endmodule

// ==== Module: i2c_master_byte_ctrl ====
module i2c_master_byte_ctrl ( clk, rst, nReset, ena, clk_cnt, start, stop, read, write, ack_in, din, cmd_ack, ack_out, dout, i2c_busy, i2c_al, scl_i, scl_o, scl_oen, sda_i, sda_o, sda_oen ); input clk; input rst; input nReset; input ena; input [15:0] clk_cnt; input start; input stop; input read; input write; input ack_in; input [7:0] din; output cmd_ack; reg cmd_ack; output ack_out; reg ack_out; output i2c_busy; output i2c_al; output [7:0] dout; input scl_i; output scl_o; output scl_oen; input sda_i; output sda_o; output sda_oen; parameter [4:0] ST_IDLE = 5'b0_0000; parameter [4:0] ST_START = 5'b0_0001; parameter [4:0] ST_READ = 5'b0_0010; parameter [4:0] ST_WRITE = 5'b0_0100; parameter [4:0] ST_ACK = 5'b0_1000; parameter [4:0] ST_STOP = 5'b1_0000; reg [3:0] core_cmd; reg core_txd; wire core_ack, core_rxd; reg [7:0] sr; reg shift, ld; wire go; reg [2:0] dcnt; wire cnt_done; i2c_master_bit_ctrl bit_controller ( .clk ( clk ), .rst ( rst ), .nReset ( nReset ), .ena ( ena ), .clk_cnt ( clk_cnt ), .cmd ( core_cmd ), .cmd_ack ( core_ack ), .busy ( i2c_busy ), .al ( i2c_al ), .din ( core_txd ), .dout ( core_rxd ), .scl_i ( scl_i ), .scl_o ( scl_o ), .scl_oen ( scl_oen ), .sda_i ( sda_i ), .sda_o ( sda_o ), .sda_oen ( sda_oen ) ); assign go = (read | write | stop) & ~cmd_ack; assign dout = sr; always @(posedge clk or negedge nReset) if (!nReset) sr <= #1 8'h0; else if (rst) sr <= #1 8'h0; else if (ld) sr <= #1 din; else if (shift) sr <= #1 {sr[6:0], core_rxd}; always @(posedge clk or negedge nReset) if (!nReset) dcnt <= #1 3'h0; else if (rst) dcnt <= #1 3'h0; else if (ld) dcnt <= #1 3'h7; else if (shift) dcnt <= #1 dcnt - 3'h1; assign cnt_done = ~(|dcnt); reg [4:0] c_state; always @(posedge clk or negedge nReset) if (!nReset) begin core_cmd <= #1 `I2C_CMD_NOP; core_txd <= #1 1'b0; shift <= #1 1'b0; ld <= #1 1'b0; cmd_ack <= #1 1'b0; c_state <= #1 ST_IDLE; ack_out <= #1 1'b0; end else if (rst | i2c_al) begin core_cmd <= #1 `I2C_CMD_NOP; core_txd <= #1 1'b0; shift <= #1 1'b0; ld <= #1 1'b0; cmd_ack <= #1 1'b0; c_state <= #1 ST_IDLE; ack_out <= #1 1'b0; end else begin core_txd <= #1 sr[7]; shift <= #1 1'b0; ld <= #1 1'b0; cmd_ack <= #1 1'b0; case (c_state) ST_IDLE: if (go) begin if (start) begin c_state <= #1 ST_START; core_cmd <= #1 `I2C_CMD_START; end else if (read) begin c_state <= #1 ST_READ; core_cmd <= #1 `I2C_CMD_READ; end else if (write) begin c_state <= #1 ST_WRITE; core_cmd <= #1 `I2C_CMD_WRITE; end else begin c_state <= #1 ST_STOP; core_cmd <= #1 `I2C_CMD_STOP; end ld <= #1 1'b1; end ST_START: if (core_ack) begin if (read) begin c_state <= #1 ST_READ; core_cmd <= #1 `I2C_CMD_READ; end else begin c_state <= #1 ST_WRITE; core_cmd <= #1 `I2C_CMD_WRITE; end ld <= #1 1'b1; end ST_WRITE: if (core_ack) if (cnt_done) begin c_state <= #1 ST_ACK; core_cmd <= #1 `I2C_CMD_READ; end else begin c_state <= #1 ST_WRITE; core_cmd <= #1 `I2C_CMD_WRITE; shift <= #1 1'b1; end ST_READ: if (core_ack) begin if (cnt_done) begin c_state <= #1 ST_ACK; core_cmd <= #1 `I2C_CMD_WRITE; end else begin c_state <= #1 ST_READ; core_cmd <= #1 `I2C_CMD_READ; end shift <= #1 1'b1; core_txd <= #1 ack_in; end ST_ACK: if (core_ack) begin if (stop) begin c_state <= #1 ST_STOP; core_cmd <= #1 `I2C_CMD_STOP; end else begin c_state <= #1 ST_IDLE; core_cmd <= #1 `I2C_CMD_NOP; cmd_ack <= #1 1'b1; end ack_out <= #1 core_rxd; core_txd <= #1 1'b1; end else core_txd <= #1 ack_in; ST_STOP: if (core_ack) begin c_state <= #1 ST_IDLE; core_cmd <= #1 `I2C_CMD_NOP; cmd_ack <= #1 1'b1; end endcase end endmodule

// ==== Module: i2c_master_bit_ctrl ====
module i2c_master_bit_ctrl ( input clk, input rst, input nReset, input ena, input [15:0] clk_cnt, input [ 3:0] cmd, output reg cmd_ack, output reg busy, output reg al, input din, output reg dout, input scl_i, output scl_o, output reg scl_oen, input sda_i, output sda_o, output reg sda_oen ); reg [ 1:0] cSCL, cSDA; reg [ 2:0] fSCL, fSDA; reg sSCL, sSDA; reg dSCL, dSDA; reg dscl_oen; reg sda_chk; reg clk_en; reg slave_wait; reg [15:0] cnt; reg [13:0] filter_cnt; reg [17:0] c_state; always @(posedge clk) dscl_oen <= #1 scl_oen; always @(posedge clk or negedge nReset) if (!nReset) slave_wait <= 1'b0; else slave_wait <= (scl_oen & ~dscl_oen & ~sSCL) | (slave_wait & ~sSCL); wire scl_sync = dSCL & ~sSCL & scl_oen; always @(posedge clk or negedge nReset) if (~nReset) begin cnt <= #1 16'h0; clk_en <= #1 1'b1; end else if (rst || ~|cnt || !ena || scl_sync) begin cnt <= #1 clk_cnt; clk_en <= #1 1'b1; end else if (slave_wait) begin cnt <= #1 cnt; clk_en <= #1 1'b0; end else begin cnt <= #1 cnt - 16'h1; clk_en <= #1 1'b0; end always @(posedge clk or negedge nReset) if (!nReset) begin cSCL <= #1 2'b00; cSDA <= #1 2'b00; end else if (rst) begin cSCL <= #1 2'b00; cSDA <= #1 2'b00; end else begin cSCL <= {cSCL[0],scl_i}; cSDA <= {cSDA[0],sda_i}; end always @(posedge clk or negedge nReset) if (!nReset ) filter_cnt <= 14'h0; else if (rst || !ena ) filter_cnt <= 14'h0; else if (~|filter_cnt) filter_cnt <= clk_cnt >> 2; else filter_cnt <= filter_cnt -1; always @(posedge clk or negedge nReset) if (!nReset) begin fSCL <= 3'b111; fSDA <= 3'b111; end else if (rst) begin fSCL <= 3'b111; fSDA <= 3'b111; end else if (~|filter_cnt) begin fSCL <= {fSCL[1:0],cSCL[1]}; fSDA <= {fSDA[1:0],cSDA[1]}; end always @(posedge clk or negedge nReset) if (~nReset) begin sSCL <= #1 1'b1; sSDA <= #1 1'b1; dSCL <= #1 1'b1; dSDA <= #1 1'b1; end else if (rst) begin sSCL <= #1 1'b1; sSDA <= #1 1'b1; dSCL <= #1 1'b1; dSDA <= #1 1'b1; end else begin sSCL <= #1 &fSCL[2:1] | &fSCL[1:0] | (fSCL[2] & fSCL[0]); sSDA <= #1 &fSDA[2:1] | &fSDA[1:0] | (fSDA[2] & fSDA[0]); dSCL <= #1 sSCL; dSDA <= #1 sSDA; end reg sta_condition; reg sto_condition; always @(posedge clk or negedge nReset) if (~nReset) begin sta_condition <= #1 1'b0; sto_condition <= #1 1'b0; end else if (rst) begin sta_condition <= #1 1'b0; sto_condition <= #1 1'b0; end else begin sta_condition <= #1 ~sSDA & dSDA & sSCL; sto_condition <= #1 sSDA & ~dSDA & sSCL; end always @(posedge clk or negedge nReset) if (!nReset) busy <= #1 1'b0; else if (rst ) busy <= #1 1'b0; else busy <= #1 (sta_condition | busy) & ~sto_condition; reg cmd_stop; always @(posedge clk or negedge nReset) if (~nReset) cmd_stop <= #1 1'b0; else if (rst) cmd_stop <= #1 1'b0; else if (clk_en) cmd_stop <= #1 cmd == `I2C_CMD_STOP; always @(posedge clk or negedge nReset) if (~nReset) al <= #1 1'b0; else if (rst) al <= #1 1'b0; else al <= #1 (sda_chk & ~sSDA & sda_oen) | (|c_state & sto_condition & ~cmd_stop); always @(posedge clk) if (sSCL & ~dSCL) dout <= #1 sSDA; parameter [17:0] idle = 18'b0_0000_0000_0000_0000; parameter [17:0] start_a = 18'b0_0000_0000_0000_0001; parameter [17:0] start_b = 18'b0_0000_0000_0000_0010; parameter [17:0] start_c = 18'b0_0000_0000_0000_0100; parameter [17:0] start_d = 18'b0_0000_0000_0000_1000; parameter [17:0] start_e = 18'b0_0000_0000_0001_0000; parameter [17:0] stop_a = 18'b0_0000_0000_0010_0000; parameter [17:0] stop_b = 18'b0_0000_0000_0100_0000; parameter [17:0] stop_c = 18'b0_0000_0000_1000_0000; parameter [17:0] stop_d = 18'b0_0000_0001_0000_0000; parameter [17:0] rd_a = 18'b0_0000_0010_0000_0000; parameter [17:0] rd_b = 18'b0_0000_0100_0000_0000; parameter [17:0] rd_c = 18'b0_0000_1000_0000_0000; parameter [17:0] rd_d = 18'b0_0001_0000_0000_0000; parameter [17:0] wr_a = 18'b0_0010_0000_0000_0000; parameter [17:0] wr_b = 18'b0_0100_0000_0000_0000; parameter [17:0] wr_c = 18'b0_1000_0000_0000_0000; parameter [17:0] wr_d = 18'b1_0000_0000_0000_0000; always @(posedge clk or negedge nReset) if (!nReset) begin c_state <= #1 idle; cmd_ack <= #1 1'b0; scl_oen <= #1 1'b1; sda_oen <= #1 1'b1; sda_chk <= #1 1'b0; end else if (rst | al) begin c_state <= #1 idle; cmd_ack <= #1 1'b0; scl_oen <= #1 1'b1; sda_oen <= #1 1'b1; sda_chk <= #1 1'b0; end else begin cmd_ack <= #1 1'b0; if (clk_en) case (c_state) idle: begin case (cmd) `I2C_CMD_START: c_state <= #1 start_a;
`I2C_CMD_STOP: c_state <= #1 stop_a;
`I2C_CMD_WRITE: c_state <= #1 wr_a;
`I2C_CMD_READ: c_state <= #1 rd_a;
default: c_state <= #1 idle; endcase scl_oen <= #1 scl_oen; sda_oen <= #1 sda_oen; sda_chk <= #1 1'b0; end start_a: begin c_state <= #1 start_b; scl_oen <= #1 scl_oen; sda_oen <= #1 1'b1; sda_chk <= #1 1'b0; end start_b: begin c_state <= #1 start_c; scl_oen <= #1 1'b1; sda_oen <= #1 1'b1; sda_chk <= #1 1'b0; end start_c: begin c_state <= #1 start_d; scl_oen <= #1 1'b1; sda_oen <= #1 1'b0; sda_chk <= #1 1'b0; end start_d: begin c_state <= #1 start_e; scl_oen <= #1 1'b1; sda_oen <= #1 1'b0; sda_chk <= #1 1'b0; end start_e: begin c_state <= #1 idle; cmd_ack <= #1 1'b1; scl_oen <= #1 1'b0; sda_oen <= #1 1'b0; sda_chk <= #1 1'b0; end stop_a: begin c_state <= #1 stop_b; scl_oen <= #1 1'b0; sda_oen <= #1 1'b0; sda_chk <= #1 1'b0; end stop_b: begin c_state <= #1 stop_c; scl_oen <= #1 1'b1; sda_oen <= #1 1'b0; sda_chk <= #1 1'b0; end stop_c: begin c_state <= #1 stop_d; scl_oen <= #1 1'b1; sda_oen <= #1 1'b0; sda_chk <= #1 1'b0; end stop_d: begin c_state <= #1 idle; cmd_ack <= #1 1'b1; scl_oen <= #1 1'b1; sda_oen <= #1 1'b1; sda_chk <= #1 1'b0; end rd_a: begin c_state <= #1 rd_b; scl_oen <= #1 1'b0; sda_oen <= #1 1'b1; sda_chk <= #1 1'b0; end rd_b: begin c_state <= #1 rd_c; scl_oen <= #1 1'b1; sda_oen <= #1 1'b1; sda_chk <= #1 1'b0; end rd_c: begin c_state <= #1 rd_d; scl_oen <= #1 1'b1; sda_oen <= #1 1'b1; sda_chk <= #1 1'b0; end rd_d: begin c_state <= #1 idle; cmd_ack <= #1 1'b1; scl_oen <= #1 1'b0; sda_oen <= #1 1'b1; sda_chk <= #1 1'b0; end wr_a: begin c_state <= #1 wr_b; scl_oen <= #1 1'b0; sda_oen <= #1 din; sda_chk <= #1 1'b0; end wr_b: begin c_state <= #1 wr_c; scl_oen <= #1 1'b1; sda_oen <= #1 din; sda_chk <= #1 1'b0; end wr_c: begin c_state <= #1 wr_d; scl_oen <= #1 1'b1; sda_oen <= #1 din; sda_chk <= #1 1'b1; end wr_d: begin c_state <= #1 idle; cmd_ack <= #1 1'b1; scl_oen <= #1 1'b0; sda_oen <= #1 din; sda_chk <= #1 1'b0; end endcase end assign scl_o = 1'b0; assign sda_o = 1'b0; endmodule
